interface pc_if(input bit clk);
   logic            rstn;
   logic            ld;
   logic [31:0]     data;
   logic [31:0]     count;
endinterface
