`ifndef MEMORY_SVH
`define MEMORY_SVH

`include "memory.sv"
`include "bram.sv"

`endif
