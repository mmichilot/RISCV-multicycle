`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:  J. Callenes
// 
// Create Date: 01/04/2019 04:49:55 PM
// Design Name: 
// Module Name: Mult4to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//  J. Callenes
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module Mult6to1(
    input [31:0] In1, In2, In3, In4, In5, In6, //32-bit inputs 
    input [3:0] Sel, //selector signal
    output logic [31:0] Out
    );

    always_comb begin
        case (Sel) //a 6->1 multiplexor
            0: Out = In1; 
            1: Out = In2; 
            2: Out = In3;
            3: Out = In4;
            4: Out = In5;
            5: Out = In6;
            default: Out = In1; 
        endcase
    end

endmodule

module Mult5to1(
    input [31:0] In1, In2, In3, In4, In5, //four 64-bit inputs 
    input [2:0] Sel, //selector signal
    output logic [31:0] Out //64-bit output
    );

    always_comb begin
        case (Sel) //a 5->1 multiplexor
            0: Out = In1; 
            1: Out = In2; 
            2: Out = In3;
            3: Out = In4;
            4: Out = In5;
            default: Out = In1; 
        endcase
    end

endmodule

module Mult4to1(
    input [31:0] In1, In2, In3, In4, //four 64-bit inputs 
    input [1:0] Sel, //selector signal
    output logic [31:0] Out //64-bit output
    );

    always_comb begin
        case (Sel) //a 4->1 multiplexor
            0: Out = In1; 
            1: Out = In2; 
            2: Out = In3;
            default: Out = In4; 
        endcase
    end

endmodule

module Mult2to1(
    input [31:0] In1, In2, //four 64-bit inputs 
    input Sel, //selector signal
    output logic [31:0] Out //64-bit output
    );

    always_comb begin
        case (Sel) //a 4->1 multiplexor
            0: Out <= In1;            
            default: Out <= In2; 
        endcase
    end

endmodule
