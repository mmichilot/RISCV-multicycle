`ifndef MEMORY_SVH
`define MEMORY_SVH

`include "sram.sv"
`include "bram.sv"

`endif
