`ifndef CPU_SVH
`define CPU_SVH

`include "cpu.sv"
`include "bus_matrix.sv"

`endif
