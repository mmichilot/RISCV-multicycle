`ifndef SYS_BUS_SVH
`define SYS_BUS_SVH

`include "sys_bus.sv"

`endif
