`ifndef SYS_BUS_SVH
`define SYS_BUS_SVH

`include "wishbone_bus.sv"

`endif
