`ifndef CORE_SVH
`define CORE_SVH

`include "alu.sv"
`include "brn_gen.sv"
`include "control_unit.sv"
`include "core.sv"
`include "datapath.sv"
`include "decoder.sv"
`include "immed_gen.sv"
`include "prog_cntr.sv"
`include "reg_file.sv"
`include "sz_ex.sv"

`endif
