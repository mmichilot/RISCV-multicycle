`ifndef SYS_BUS_SVH
`define SYS_BUS_SVH

`include "otter_bus.sv"

`endif
